LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE UC_pack IS

	TYPE states_UC IS (INICIO, INICIO_PARTIDA, PARTIDA, GAME_OVER);

END PACKAGE;
